module terminate(
    input a
    );


endmodule
