module calculator(
    input a
    );


endmodule
